`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   00:16:11 08/27/2025
// Design Name:   Dual_Core_Top_io_sim
// Module Name:   D:/Ido_Matan/Project_A/HOME_VER/Dual_Test.v
// Project Name:  HOME_VER
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: Dual_Core_Top_io_sim
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module Dual_Test;

	// Inputs
	reg CLK_IN;
	reg RST;
	reg PC_step_en;

	// Outputs
	wire AS_N;
	wire WR_N;
	wire [31:0] AO;
	wire [31:0] DO;
	wire PA_success;
	wire PB_success;
	wire PA_pass;
	wire PB_pass;
	wire in_idle;

	// Instantiate the Unit Under Test (UUT)
	Dual_Core_Top_io_sim uut (
		.CLK_IN(CLK_IN), 
		.RST(RST), 
		.PC_step_en(PC_step_en), 
		.AS_N(AS_N), 
		.WR_N(WR_N), 
		.AO(AO), 
		.DO(DO), 
		.PA_success(PA_success), 
		.PB_success(PB_success), 
		.PA_pass(PA_pass), 
		.PB_pass(PB_pass), 
		.in_idle(in_idle)
	);

	initial 
	 CLK_IN = 1 ;
	 always #50 CLK_IN = ~ CLK_IN ; 

	initial begin
		// Initialize Inputs
		RST = 1;
		PC_step_en = 0;

		// Wait 104 ns for global reset to finish
		#104;
		
		RST = 0 ;
		
		
		
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		
	
	
	
	
			PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
			PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		
		
		
		
		
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;
		PC_step_en = 1;
		#100;
		PC_step_en = 0;
		#1500;



	end
      
endmodule

